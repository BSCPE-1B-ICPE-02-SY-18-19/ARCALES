CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 110 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
77070354 0
0
6 Title:
5 Name:
0
0
0
11
6 74LS48
188 959 485 0 14 29
0 3 4 5 6 26 27 9 10 11
12 13 14 15 28
0
0 0 4832 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5130 0 0
2
43529.9 10
0
6 74112~
219 292 499 0 7 32
0 7 7 8 7 7 25 6
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
391 0 0
2
43529.9 9
0
6 74112~
219 439 499 0 7 32
0 7 6 8 6 7 24 5
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3124 0 0
2
43529.9 8
0
6 74112~
219 608 496 0 7 32
0 7 16 8 16 7 23 4
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3421 0 0
2
43529.9 7
0
6 74112~
219 755 498 0 7 32
0 7 17 8 17 7 22 3
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8157 0 0
2
43529.9 6
0
9 2-In AND~
219 515 363 0 3 22
0 6 5 16
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
43529.9 5
0
9 2-In AND~
219 683 371 0 3 22
0 16 4 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
43529.9 4
0
9 CC 7-Seg~
183 894 264 0 17 19
10 15 14 13 12 11 10 9 21 2
0 0 0 1 1 1 1 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7361 0 0
2
43529.9 3
0
7 Pulser~
4 91 469 0 10 12
0 18 19 8 20 0 0 5 5 5
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4747 0 0
2
43529.9 2
0
2 +V
167 292 419 0 1 3
0 7
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
43529.9 1
0
7 Ground~
168 978 151 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
43529.9 0
0
37
1 9 2 0 0 0 0 11 8 0 0 4
978 159
978 201
894 201
894 222
0 1 3 0 0 0 0 0 1 7 0 5
796 462
796 607
892 607
892 449
927 449
0 2 4 0 0 0 0 0 1 29 0 5
639 460
639 615
900 615
900 458
927 458
0 3 5 0 0 0 0 0 1 27 0 5
481 463
481 621
906 621
906 467
927 467
0 4 6 0 0 0 0 0 1 37 0 5
331 463
331 630
913 630
913 476
927 476
0 1 7 0 0 0 0 0 10 24 0 5
236 463
235 463
235 436
292 436
292 428
7 0 3 0 0 0 0 5 0 0 0 2
779 462
809 462
1 0 7 0 0 0 0 10 0 0 12 2
292 428
292 428
0 0 7 0 0 0 0 0 0 12 15 2
353 428
353 526
1 1 7 0 0 0 0 4 5 0 0 4
608 433
608 428
755 428
755 435
1 1 7 0 0 0 0 3 4 0 0 4
439 436
439 428
608 428
608 433
1 1 7 0 0 0 0 2 3 0 0 4
292 436
292 428
439 428
439 436
5 5 7 0 0 0 0 4 5 0 0 4
608 508
608 527
755 527
755 510
5 5 7 0 0 0 0 3 4 0 0 4
439 511
439 527
608 527
608 508
5 5 7 0 0 0 0 2 3 0 0 4
292 511
292 526
439 526
439 511
3 0 8 0 0 0 0 9 0 0 34 4
115 460
138 460
138 561
211 561
7 7 9 0 0 0 0 1 8 0 0 5
991 449
1023 449
1023 337
909 337
909 300
8 6 10 0 0 0 0 1 8 0 0 5
991 458
1018 458
1018 332
903 332
903 300
9 5 11 0 0 0 0 1 8 0 0 5
991 467
1013 467
1013 327
897 327
897 300
10 4 12 0 0 0 0 1 8 0 0 5
991 476
1008 476
1008 322
891 322
891 300
11 3 13 0 0 0 0 1 8 0 0 5
991 485
1003 485
1003 317
885 317
885 300
12 2 14 0 0 0 0 1 8 0 0 5
991 494
998 494
998 312
879 312
879 300
13 1 15 0 0 0 0 1 8 0 0 5
991 503
993 503
993 307
873 307
873 300
4 2 7 0 0 0 0 2 2 0 0 4
268 481
236 481
236 463
268 463
2 0 16 0 0 0 0 4 0 0 26 2
584 460
546 460
0 4 16 0 0 0 0 0 4 28 0 3
546 363
546 478
584 478
2 7 5 0 0 0 0 6 3 0 0 4
491 372
490 372
490 463
463 463
3 1 16 0 0 0 0 6 7 0 0 4
536 363
546 363
546 362
659 362
2 7 4 0 0 0 0 7 4 0 0 4
659 380
650 380
650 460
632 460
2 0 17 0 0 0 0 5 0 0 31 2
731 462
710 462
3 4 17 0 0 0 0 7 5 0 0 4
704 371
710 371
710 480
731 480
3 0 8 0 0 0 0 4 0 0 34 3
578 469
565 469
565 562
3 0 8 0 0 0 0 3 0 0 34 3
409 472
393 472
393 562
3 3 8 0 0 0 0 2 5 0 0 6
262 472
211 472
211 562
700 562
700 471
725 471
1 0 6 0 0 0 0 6 0 0 36 3
491 354
373 354
373 463
4 0 6 0 0 16 0 3 0 0 37 3
415 481
373 481
373 463
7 2 6 0 0 0 0 2 3 0 0 2
316 463
415 463
2
-37 0 0 0 400 255 0 0 0 3 2 1 49
8 Consolas
0 0 0 35
150 122 863 183
169 131 843 174
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
-29 0 0 0 400 0 0 0 0 3 2 1 49
8 Consolas
0 0 0 17
14 29 298 77
28 36 283 70
17 ARCALES, KLIEN T.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
